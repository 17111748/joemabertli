`define A_N        1
`define A_M        3
`define B_N        3
`define B_M        1
`define TEST_CASES 1
`define BITWIDTH   4
`define TIME_MAX   2147483647

`define FAIL_ON_ERROR
