`define A_N        16
`define A_M        16
`define B_N        16
`define B_M        16
`define TEST_CASES 1
`define BITWIDTH   4
`define TIME_MAX   50000

// `define FAIL_ON_ERROR
