/*
`define A_N          2
`define A_M          2
`define B_N          2
`define B_M          2
*/
`define DIM          2
`define BITWIDTH     8
`define OUT_BITWIDTH 16
`define TIME_MAX     1000000
`define MAX_TRACES   10

`define FAIL_ON_ERROR
