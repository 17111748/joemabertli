
`define DIM          8

`define A_N          8
`define A_M          8
`define B_N          8
`define B_M          8

`define BITWIDTH     8
`define OUT_BITWIDTH 16
`define TIME_MAX     1000000
`define MAX_TRACES   1
`define TEST_CASES   1

`define FAIL_ON_ERROR
