`define DIM 8
`define BITWIDTH 8
`define OUT_BITWIDTH 16
`define TIME_MAX 30000
`define MAX_TRACES 3
`define FAIL_ON_ERROR