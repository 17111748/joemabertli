`define A_N        4
`define A_M        4
`define B_N        4
`define B_M        4
`define TEST_CASES 1
`define BITWIDTH   4
`define TIME_MAX   50000

`define FAIL_ON_ERROR
