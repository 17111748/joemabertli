`define DIM          2
`define BITWIDTH     8
`define OUT_BITWIDTH 16
`define TIME_MAX     1000
`define MAX_TRACES   10

`define FAIL_ON_ERROR
